----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:28:47 10/02/2020 
-- Design Name: 
-- Module Name:    LED - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity LED is
    Port ( DPSwitch : in  STD_LOGIC_VECTOR (4 downto 0);
           SevenSegment : out  STD_LOGIC_VECTOR (7 downto 0);
           Enable : out  STD_LOGIC_VECTOR (2 downto 0));
end LED;

architecture Behavioral of LED is

begin


end Behavioral;

